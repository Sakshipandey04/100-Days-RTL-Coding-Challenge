`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Create Date: 22.08.2025 19:29:27 
// Module Name: sr_ff ///

module sr_ff(
   input S, R,
   input clk,
   output reg Q
    );
    
    initial Q=0;
    always@(posedge clk)begin
    case({S,R})
      2'b00: Q <= Q;
      2'b01: Q <= 0;
      2'b10: Q <= 1;
      2'b11: Q <= 1'bx;
    endcase
  end
      
endmodule
